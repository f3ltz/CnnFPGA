module lenet_TB ();

reg [32*32*16-1:0] input_ANN; 

reg clk, reset;
wire [3:0] output_ANN;
reg [5*5*6*16-1:0] Conv1F;
reg [400-1:0] memory1 [0:6-1];
reg [5*5*6*16*16-1:0] Conv2F;
reg [5*5*6*16-1:0] memory2 [0:16-1];

integer i;
integer code;
integer fd ;

localparam PERIOD = 100;

always
	#(PERIOD/2) clk = ~clk;

initial begin
  
    #0
    clk = 1'b0;
    reset = 1'b1;
//     label:3
//    input_ANN = 16384'h3413345332253125341335133326341334933413332634133413322531a530a5322534133493345334d335d33593361335d3375437d437d437d4384a390a39ea3493355333a631a533a63413322533a632a634d334d334533326312531a532a63326349334d334533553369336d4375435d3369336d437d437d4386a392a398a351335933493332635133326322532253326332633a634933413332633263326322533a6351338aa396a3aca3aca39aa396a380a369337d43794380a388a396a3553351335133225341331a530a530a532a632252e4ab4afa9703493332632a633a634933a8a39ca398a39aa3b8b3c653bcb3c5539ca382a37143754380a38ca355334133326322532a633a630a5322533a632a62523bd2cb6af345334d335533a2a3cd53beb3794361335d3384a392a3beb3b0b3bab3a4a386a3754388a38ca355336d437d434d3332633a6322532a6345332a63225b0dd302537943b2b3d263cb53cd53a6a3553332633263513390a388a39aa3ce53cd53a0a365337d4386a380a38ca3e163bcb33a6312532a6312531a532a631a53593380a365339ca3c553aeb3bcb3a8a2d49aeb93413386a380a36133a8a3c353d963c7537d43754388a349338ea3dd63c853553322533a63225302533a635d338ca35d32a9236d43a2a394a3a2a3b6b3413b4ef30a5392a388a392a3aca3cd53d463d763a2a36d4382ab6af37d43ce533262f4a341332a630252f4aaeb9394a36d4b05db0dd35933aca3aca3a6a3b2b3bcb3025a6e037943aeb3b2b3a8a3beb3cf53e363ca536933714b918a970388ab46fb42f332633a632a6ba18bd3cba58a6e0b5af1c8835533a0a3a6a3bab3ce53c2530251c8830a5388a3aaa3a4a3a6a3b8b3d663e863b4b3754b9d83553b2ddb818b5af34533225392abc0cbdcdbbf9afb9b7b0aeb9359335933b6b3aeb3db63a2ab7f0b2ddb25d384a3a6a382a3a0a3b2b3cc53e263d763a6abad83714aeb9b8d8b83830252d49386a386aba58b978b2ddb7f0b8f832a6369338aa3a8a3e163326bc3cb46facb839ca3aeb394a380a3a2a3b8b3d153cf53cc5bb39390a2892b978b5ef2d492c4934933babb5afb2dd3413b858bc4cb35d3553351335533d56b1ddba98b35d341339ea3a8a3a6a392a3a2a3a2a3bcb3bab3ce5baf8390ab4afba98361336532c4931a53b2b1c882f4ab42fb918bd1cb8b82a92341335533c05b42fb9d8b0dd36133a4a3aeb3beb3b0b388a386a39ea39ca3b8bbb7936d4b818ba5836d439ca31a52f4a3b4b37143125ba78b9d8b7b0adb9b0dda970386a3c05b42fb91825232f4a36933a4a396a390a36933513390a3a4a38eabbb92c49b838b9981c883aca32a62f4a390a33a62892bd7dbe5dacb82c493225359337d439ca1c88b62fb1dd36d43a4a3c0539ea37d4369336133a0a38aa3714bc3cb25db7f0ba38b8583a6a31252f4a32a63aebb0ddb770b4af289237543754386a384a394ab1ddacb8adb92d4937943b6b3b0b394a394a3a0a392a35133693bcfcb7f0b818ba38b9b8386a38cab3dea6e0394a341336d437d43754396a365339ca384a2d49388a3ce5332630253c153ce53cf53c15392a38ca34d333a63593bcbcb9f8b8d8b998b9d82e4a39eaacb8b2dd2f4a394a3c45322535933413afb939aa392aacb834133693386a3c253cb53dd63c853c0536d4322531a5341334d3bb39ba98b8f8b958b9b8b25d39aa32a631a5a1bea1be3ca533a6388aa1beb93834933bab332630a52e4a3a2a3d663d463d6639aa38ea30a52e4a332634533593b5afbb39b958b8d8b9b8b52f380a1c88b8f83794398a3b4b39aa3413b8d8ba18b2dd386a3aeb3b2b3cb53d563db63e863d053c25386a30a531a5369335d3379433a6bbf9b938b898b998afb93a2ab46fbefdbd5da970acb8b4efb9b8bb99bb39b8982a9236933c953d963d563c553b4b3aca3b0b394a392a38aa39aa3a6a3aaa386abb18b9b8b8d8b958b0dd3613bcbcbf4dbf5dbd4cab712e4aa9702c492a92332639ea3a8a3b2b3b2b3b4b3b2b3a2a3a0a3a8a3a4a396a38ca3a2a3a4a3a8a3aeb2f4ab6efb8d8b9d8b838b770becdbf2dbddd2d493aaa3b8b3c053c053c353bcb3bab3bab3bab3b6b3aca3aeb3b0b3aeb3a6a3a4a3a0a39ea3a2a3a0a3aca3b2b3b8b394ab2ddb9181c88bad8bf2dbecdb4ef39ea3b2b3b2b3b0b3b4b3b4b3b2b3b8b3bcb3c253bcb3b6b3b6b3aeb3a8a392a390a394a394a39ca3a4a394a38aa3aeb3bab386ab05d2523bcdcbf5dbb9939ea3a6a3aca3a8a3a8a3b6b3b8b3bab3bcb3c053bab3b6b3b0b3aaa3a4a38aa386a386a38aa38ca392a35d330a5384a3a4a3b8b3b8b39aaaeb9bdcdbecda9703a6a3aeb3a0a3a4a3b8b3b8b3b6b3b4b3b8b3b4b3b0b3aca3a2a390a388a390a3a0a3a4a3aeb38ca34533025351338aa3a4a3b4b3b6b3b6b384abd0cbd8d3413390a3a2a3aeb39ca3b0b3beb3b8b3b4b3aeb3aca3aca39ea3aca3aaa398a39aa3aaa3bcb39ca349335533a0a3a0a38ca3a6a3aeb3b2b3aeb3b4b3025baf8398a3a0a3a4a3a2a390a398a3a0a3b6b3beb3bcb3aeb3a6a3a8a3a6a3aaa3aca3b0b3aaa39aa359338ca3b2b3d463a4a359339ea3b4b3aca3b2b3aeb3beb388a3aeb3c553c953bcb3a6a398a394a3a6a3a0a396a398a39ca3a2a3a6a3b2b3bcb3aca382a32a6341337d43a4a3d153b6b3794398a3b8b3a8a3aeb3aaa3b0b3beb3b6b3c953cd53c653c953c753c053b2b3a0a394a386a365337d43a2a3b0b3b0b38ea3326b1dd1c8837d43c053c053cf538ca390a3aca3b0b3b0b3aca3b4b3beb3c153cb53ce53c753cb53c753d153d563c953b0b390a3693384a3a0a3a2a3b0b384a3225a97030a539ca3c453bab3cd5;
    // label:8
//    input_ANN = 16384'hbe3dbdfdbe0dbe0dbe0dbe0dbe0dbe0dbe0dbe0dbe1dbe1dbe1dbe1dbe1dbe0dbe0dbe0dbe0dbe0dbe0dbe0dbe0dbe1dbe0dbe1dbe0dbe0dbe0dbe1dbe1dbe0dbe6dbe3dbe3dbe3dbe3dbe3dbe3dbe3dbe3dbe3dbe4dbe4dbe4dbe4dbe4dbe4dbe3dbe2dbe4dbe3dbe3dbe2dbe4dbe4dbe4dbe4dbe3dbe3dbe3dbe4dbe4dbe3dbe5dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe2dbe3dbe2dbe2dbe2dbe3dbe3dbdddbe2dbe1dbe2dbe2dbe2dbe2dbe2dbe2dbe3dbe3dbe2dbe6dbe3dbe3dbe3dbe3dbe3dbe3dbe3dbe2dbe2dbe2dbe2dbe2dbe2dbe3dbe3dbe1dbe0dbdedbdadbaf8bcecbc9cbdcdbe3dbe2dbe2dbe2dbe2dbe3dbe3dbe3dbe5dbe2dbe3dbe3dbe3dbe3dbe3dbe3dbe2dbe2dbe3dbe3dbe2dbe2dbe3dbe3dbe5dbe4dbd8dbc9cb858bc2cbd1cbdedbe4dbe3dbe3dbe3dbe4dbe4dbe4dbe4dbe7dbe3dbe3dbe3dbe3dbe3dbe4dbe3dbe2dbe3dbe4dbe4dbe3dbe1dbe4dbdfdbcecbc2cbb79ba38b918bb39bcdcbdcdbe4dbe4dbe4dbe4dbe4dbe5dbe5dbe5dbdddbdbdbdfdbdddbe1dbe4dbe5dbe4dbe4dbe4dbe5dbe6dbdcdbdbdbe4dbd9dbb59b8f8b8f8b878b5efb52fb7b0bc4cbe5dbe4dbe3dbe3dbe4dbe5dbe5dbe6dbd2cbdddbe1dbdfdbe1dbe4dbe5dbe5dbe6dbe6dbe5dbe7dbc3cbd5dbe3dbd1cbc1cbbb9bbb9ba78b978b878b8b8bb99be4dbe5dbe4dbe5dbe5dbe6dbe6dbe6dbdddbe0dbe3dbe3dbe4dbe4dbe4dbe4dbe5dbe5dbe5dbe7dbbb9bd4cbe1dbdedbcccbcfcbdadbd0cbd3cbd5dbdddbdfdbe4dbe3dbe4dbe5dbe5dbe6dbe7dbe6d25232892a970b35dba18bdfdbe3dbe3dbe2dbe3dbe4dbe4dbcfcbdbdbe1dbe5dbdedbdedbe3dbdfdbe3dbdddbcecbbf9ba38b918b938bb79bdfdbe7dbe7dbe7d3125349333263225b52fbdbdbdbdbdbdbe1dbe2dbe2dbe3dbe1dbe2dbe4dbe2dbe3dbe4dbe3dbdedbc2cb978b62fb3deb15da9702c49b5efbd9dbe7dbe6dbe7dbc8cbbf9bc9cbc9cbd0cbdadbcdcbc9cbcecbd5dbd8dbd1cbd0cbd2cbd7dbdbdbe0dbe1dbe2dbdcdbbd9bb18bb79bad8bb79b958b35dbb39bdbdbe5dbe7dbe7dbc5cbc0cbcacbd2cbdadbd2cbc7cb8b8b978bcbcb9b83693369334d331252523b2ddb72fbcccbe0dbdcdbdedbdfdbd8dbdbdbd2cbc2cbdcdbd9dbdcdbe5dbe7d3025322532252c49b0ddb998bbd9bbb9bd1cbdadb8383c353c653c353c253aeb35d3b7f0bdadbe6dbe4dbdedbdbdbcacbc7cbd0cbd1cbc5cba38bb79bd3cbdcd3b2b3a6a3b4b3aaaa6e0b3deb52fbbf9bd8dbd2cb918345336933553b2ddbad8bcccbd7dbd4cbc5cba58b770b46fa6e02c49a6e0b05dacb81c88b2ddbb39bc8c3d363c2538eaacb8b15d37d43493b62fb958baf8baf8bad8bb18bc7cbdadbc8cb978b72fb35da1be31a536d437d43693351334532a92b25db66fb858bc1cbbd93f663e96ab71bcdcb15d32a6a1beb770b9b8bc9cbd7dbe0dbdfdbe6dbe2dba38b4efb35db4efb5efb818b6afb6afb818b878b8d8ba78bc0cbc3cbb18b978b87840033c85bc6cbdfdbc3cbc5cbcdcbd9dbdedbe4dbe5dbe4dbd1cbe2dbe1dbd7dbcdcbb99bcbcbc7cbc7cbcacbc8cbc0cbab8ba78b938b62fb42fafb9acb8b35d3d96b4efbc2cbb79bb79bc7cbc8cbc6cbc5cbc2cbc5cbc4cbad8bb79b878b770b5efb838b66f2d492892b42fb0dd2d49361336d43653361333262c49ab71acb82523b938b5efb46fb35db2ddb25db2ddb2ddb15db15db25db1ddafb931a5341334532892302536933613355336d4384a38ea384a3693351333a631a52c49adb93a4a39ea39aa394a38aa382a380a37543613341331a52d491c88a1be2892252325232d49312534933693384a38ea396a392a38ca38ca38ea380a34132892b15d3f063fd63f763ed63ec63ec63ec63e863e363dc63d463cc53c353b6b3b0b3aaa3a0a39ea3aca3bcb3c353c353c353c253c053b8b3a0a38aa35d331a51c88b05d3db63f863fb63de63db63ed63fb63ff640133b0b3b0b3aca3f963f563f563f263ea63e063e563e663e263de63d763cf53c15396a3493312534d33225a6e0b5af3df63ec63f663e263b2b3c053d563e963f76400b4023bdcd3f463c653d763e863ed63ed63ec63e663de63d153beb38ca30a5a6e03125369335932892b35db9183f763fc63ff63fe63da63cf53d863e563f56401b402b3b4b3ff63413b66f2c49355337143754369335d331a5a1be1c883593396a38aa34932d49b0ddb838baf83e063fd63b0b3b0b3ff63f563f463f96400b402b4033402bbdbd3c95b15db4afb35db15db05da6e02d49359339aa3b4b3b2b38ea34132d49a970b5efb958bb393bcb3ec6403340333e8640133ff64013402bb998b998b42f40333f563b0b38ea394a394a398a3aaa3c553d153cd53aca3613312530a52a92b35db878b9d8bb5939ca3d6640334033b998402b4023b42fb998b998b998b9983e863fd63ca53a2a3b0b3c153d053d963d463c05392a355331a531a531a5a1beb46fb8d8ba58bb9938aa3ce5400b402b3e86402b402b402b4033b998b99840333b0b3e563da63c153d763e863e463c95396a35933225322532a630252a92adb9b4efb878ba78bbd9392a3d863f363fc63ff63ff64003401340234023402340233aca401b3f163e363e463d463b6b384a3493302531a5332631a51c88b05db35db72fb978bb18bbd939aa3d463e063e763ec63ee63f163f363f463f463f363f263ef63ec63e163ce53b8b396a37d4355331253225341332a62f4a1c88b0ddb4efb7f0ba18bb79bbb9392a3c353ca53cf53d363d663d663d463d463d263d053cd53c953c453aeb38ea379435d3341333a6312533a633a630252a92adb9b1ddb56fb7b0b958bad8bb99;
    // label:0
//    input_ANN = 16384'hb4efb8f8b998bb39ba38b878b898b898b8d8b998ba38ba58ba58ba58b9f8b9f8b9b8b998ba18ba58ba78ba78ba98bab8ba78ba78ba98bb79bbf9bbf9bc3cba18b4efb938ba18bb99baf8b6efb62fb72fb72fb818b8b8b958b898b8f8b770b818b8b8b7f0b838b818b858b918b898b878b898b918bb39bc6cbc7cbc8cbcdcbab8b4afb8f8b9f8bb79bc0cbad8b978b918b838b958bab8bb99bb99bbd9baf8bab8bbb9bb99bb79bb99bbb9bbf9bb79bb39bb59bbd9bc7cbc8cbc8cbc8cbcdcbad8b4afb8f8ba18bb39bbd9bb99bb39b2dd2c49b818b878b858b918b770b770b7f0b998b938b978b9f8b9d8b998b9d8b8b8bb99bc7cbc6cbc6cbc8cbc8cbcccbab8b4efb8d8b9f8bab8bb79bb79bb18b2ddb1ddb56f2a922892adb9acb8ab71aeb9b0ddadb9aeb9b1ddafb9adb9b46fa1beb8f8bc5cbc3cbc4cbc8cbc6cbcdcbaf8b42fb898b9f8ba98bb18bb59bad8b6efb978b918b5efb898b918b62fb6efb838ba18ba38b9b8bb39b9d8b9f8bad8b9f8bc1cbc9cbc8cbcacbcbcbcbcbd0cbb18b42fb838b9b8ba98bab8bb39b7f03025b6afb72fb5efb7b0b6afb0ddb3deb5afb858b7b0b9b8b938b7f0b9b8b7f0b938b838b958bc4cbc7cbc8cbc8cbcdcbad8b52fb858b958ba58bad8ba58b15d2523b15db3deb3deb05db66fb42fb3deb35db2ddb15db42fb35da1beb4afb1ddb8b8aeb9b35dbb99bc2cbc3cbc2cbc8cba78b6efb8d8b938ba38bad8ba38b8f8b9d8b858b858b8f8b878b978b8b8b8d8b918b978b998b9b8b998b838b958b998bad8b9d8ba18bbd9bc2cbc1cbc1cbc7cba38b8b8b9d8b938ba38ba78ba98bb39ba18b66fb770b66fb72fb5efb56fb6efb72fb858b8d8b898b6efb66fb770b72fb978bc3cbc1cbc0cbc2cbc3cbc2cbc6cb9f8b958bb59b9d8bab8bab8bad8bb18b9f8b6efb7f0b770b5efb72fb7f0b878b8d8b878b818b7b0b858b7f0b8b8b898b978bc0cbc0cbc0cbc0cbc1cbc0cbc6cba18b9f8bc1cbaf8bbf9bbd9ba18ba98bb99bb18baf8bb18bb18bb39bb79bbf9bbf9bbf9bbb9bb99bb99bb79bb79bbb9bbd9bbf9bc0cbc0cbbf9bc0cbbf9bc7cba78ba38bc2cbb99b978b72facb8b4efbbb9bc4cbc1cbbd9bbb9bbd9bc0cbc2cbc3cbc2cbbf9bbd9bb99bb99bbd9bbf9bbd9bbf9bc1cbc3cbc5cbc7cbc7cbcccbad8ba58bc6cbbd9b7b0aeb932a6390a3693b0ddb9b8bc0cbc0cbbd9bbf9bc2cbc5cbc5cbc5cbc6cbc4cbc2cbc2cbc5cbc5cbc4cbc3cbc3cbc3cbc3cbc3cbc6cba18ba58bc9cbc6cbc6cbc4cbaf8afb9398a3aaa380ab05db9f8bbf9bc5cbc8cbc8cbc8cbc8cbc8cbc3cbbd9bbd9bbf9bbb9bbb9bbb9bbb9bbb9bbb9bbb9bc3cb9b8ba18bcbcbc8cbc7cbc7cbcacbc6cb95834d33a6a392a2d49b918bc5cbcbcbc8cbc6cbc3cbc3cbc2cbbf9bc0cbc2cbc1cbc0cbc2cbc1cbbf9bbd9bbd9bc2cb998ba58bcdcbcccbcecbcdcbcdcbcccbd1cb918396a3b8b39ea380aacb8b9d8bc5cbc9cbc5cbc1cbbf9bbf9bc1cbc1cbc0cbc0cbc2cbc1cbc0cbc1cbbf9bc2cb9d8ba78bcecbcecbd2cbd2cbd1cbcecbcbcbc5c31a53c253a8a3aeb3aaa38aa2c49b7f0bad8bc3cbc4cbbd9bb79bc1cbc0cbbf9bc0cbc0cbbf9bc1cbbf9bc3cb9f8bab8bd0cbcccbd0cbd0cbd0cbcecbcbcbcdca6e03c053a6a3b0b3aca3aaa3b0b3a4a380a2f4ab46fb6afb9d8bc4cbc7cbc5cbc2cbc0cbbd9bbf9bbd9bc1cb9b8ba98bd1cbcdcbcfcbcfcbd0cbcfcbd0cbc5c35933d963cf53cb53c053aeb3a4a3a8a3b4b3c153c953cc53aeb31a5b62fb9b8bb99bc5cbc6cbc4cbc1cbc3cb9d8ba98bcfcbcacbcbcbcccbcfcbcdcbcdcb52f38ca3cb53e463d663c753c353aeb3a4a3a6a3a6a3beb3cf53d863c853c053b2b37142892b5efba18bb99bc3cba38ba18bc9cbc7cbc9cbcacbcbcbcdcbc1cb1dda1beb15d388a3d963d363d76396ab42fb5ef2f4a3beb38aa35d339ca3c553c452c49b7b0b6efb878b9f8bb99b958b9f8bc9cbc6cbcacbcccbcccbcdcbcbcbcbcbcbcbcfcbb18b25db25db2ddb818bc2cbc9cbb79b56fb7b0b9b8b998b6afb5efb9b8bb59bbd9bbd9bb79bbb9b958b8d8bb79bb99bb99bb79baf8ba98ba58ba38b9d8b9f8b998b938b918b8f8b918b8b8b7b0b818b8d8b898b818b898b958b938b7f0b5efb5afb6afb7f0b8f8b62f361337143593371437d4386a38ca38ea396a39ca394a3a2a3a6a3a6a39ea379434533513359335533513349334133326312530252f4a302530a530252892302534533513351334d334d3355334d334d335933513359335d335d3361335d33653345334d33693361335d33653379436d43653361335933593380a388a388a386a3553382a37143693369337d4388a392a390a394a39ea3a2a3a8a3b0b3aeb3b0b3aca3b0b3c053c353c453c653c653c753c753c653c653c753ca53ce53c6539aa3a8a3cd53c653c653c753c753c953cb53c653c853cc53d053cf53cc53cb53c953c953c653c853ce53d053cf53cd53cc53cd53cf53cf53cf53d153c75380a35133a6a3cb53c753c753c753c653ca53c853c453c953cb53cd53cd53cd53cb53cb53c753c653ca53cc53cd53ce53cc53cd53ce53ce53cc53ca53aca33263225398a3aeb3d153ca53ce53cf53cc53ce53cc53cb53cd53cf53d153cb53ca53cc53ca53c653ca53cd53ce53cb53ca53c953ca53c953cb53c5538ea30a536d43c053c253aaa3cd53c753c853c953c953c953c953c953ca53c753b0b3aeb3b4b3b8b3b4b3a6a3aca3aca3b0b3b4b3c753c953c853cb53b8b36132f4a394a3c953c953c253aca3d153cd53ce53cc53cb53ca53cc53cb53cb53cc53c253c053c053c253c353c053c053bcb3bcb3bcb3c953c953c653aeb359335933b0b3c953ca53c853c45;
    // label:6
//    input_ANN = 16384'h3c653b6b3ce53e063ea63d563c853c453c253cc53f763ed63cb53c653c953cc53b4b37543653371435d338ca3bab3c0531a533a63d563aeb3a0a3cc53c453b0b3bab394a3c353df63d663aeb3c053c053bab3d363fa63e063aeb3aaa3c353c85392a380a38aa392a37d438ca3c453bcbacb82e4a3e163ce53c753cb53aeb3bcb3a2a388a3aca3d663bab396a3beb3b6b3b2b3da63f763d563b6b3b0b3cd53d46398a39aa3c253bab384a382a3cd53b6bb25d28923ea63d663b4b39ca39ea3d05379439aa396a3c7538ea39ea3b6b3a6a3aca3e163f163d763cf53ca53d763d8638ea36d43a0a3a2a37d4384a3ca53acab35dadb93cf53a4a361335933aaa3da6365338ca33a63aca386a3aca3b0b3a6a3aca3e763f263e963df63d863c753b6b398a38aa394a39ca396a38ca3c75394ab4afb6af384a37d434d33493398a388a38ea394a398a39ea3a6a3b4b3aca3c153b4b3ea63f163e363c653aeb396a394a39ca39ea3a0a3c253d5638aa3a2a396ab62fb938349335d335532d49322536133a6a3a8a3de63c153aca39aa3a4a3ce53c753ef63e563b2b3714365336133a6a3d763c8537143d463e763653386a392ab8d8ba38302530a53125b25d392a3d153b8b3beb3e26398a394a39ea39ea3c453d563f763c75341334d3349338ea3e563f363cf537943c053d15355337943326b66fba58a6e0a9701c88b05d3cd53ef63a2a3c553c753125a6e037d43beb3a2a3c453e06388a3225351335133d263f563ca536533aaa3b0b36d430252523aeb9b4afb7f0a970acb8a6e02a923e263f16384a3c153c252523b2ddaeb93b6b3c853b2b3a4a31252f4a32253aaa3ec63d86365330a5384a35931c88ab71a6e035d3b4afb66facb8afb9a6e036133f463ef637543c153c652a92b35db42f34d33cd53d86384a312534533225398a3c5538ca341334d33025a9701c88b1dd382a3babb5afb6afab71b05d289237543f763f1634d33c953cc530a5b1ddb46fb3de3a2a3c65341334d3371434d3380a2a92b4afafb9a970289230a5345332a637943453b8d8b4ef2892b15da6e036533f663fd6384a3d463d2636933225b2ddb52fa97028921c88341333a63225390a384a2892acb825232f4a341331a536d4349330a5b6efb5ef33a62d49b1dd37143f163de636d43b4b3c15379434d32f4ab56fb56fb25d30a5289231a5322533a6351335d33693365332a62d491c8830a51c8833a6adb9b3de2f4aa6e0b3de380a3cc539ca33263a2a39ca365334133794b42fb4afa9703593369334d32f4a2a92b05d1c8830a531a535d334d333a63225b15db25db15d3326a6e0aeb9adb937943c553a2a36533aeb3aaa371434d33593ab71b42fb25db8f831a53c1536532f4a3025afb9b62fb2dd2a9231a530a537542523b838b72fb05d3125b0dd25233c253ea6392a382a398a39ca36132e4aab71a6e0b2dd2e4ab7f0b8983bab382aa970b05db15d2523adb9b72fb6afb7f0b4ef2e4a2e4ab878b9b8312525232e4a3d153d962e4a380a382a34133513252335532c4931a52c493326b898b52f30a52892b42fb42fb1ddb05da6e0afb9acb8b1ddb4efa970b25d2892b3de349332a639ca3d46380a35d33693a6e028922e4a39ea35d337542c49345332a6baf8b35d34d3aeb91c88b62fb7b0b42fb5efb56fa970b35db25dab7130a538ca3aeb392a37543a2a3125312531a5ab7137d4369339aa3a6a35533225aeb9398a2f4ab8b8adb9b3deb770b4efb46fb878b878b0dd2523b1ddb1dda1be25233bcb3a2a3b8b3b6b2523b52fa1be3025380a3a2a36d439aa3bab3413398a37542e4a3c253413b7b0b5efb8d8b858b4afb6efb8b8b35daeb9b42fb2dd2c4930a53754379439ea3693ab71aeb9adb936933c653513345339aa39ea365336933aebacb8355339aab3deb9f8b8b8b7f0b958b35db25db2ddadb92523afb92e4a322535d3394a3413b56fa1be2a9230a5390a3b8b359331a537543a2a380aa1be2f4a37d4a97030a5b25db8d8b9f8b858b898b6efb0dd2c49b05db0ddb15dadb925233493380aacb8b05d2f4a2f4a3513382ab05db9f8b62facb837d438ca2e4aadb937d438eab0ddb6efb56fb958b7f0b5efb62fb0ddaeb9b46faeb9b35dafb9252333262d49ab7130251c882f4aa1beb4afbb59bcccbbf9b878b2dd2e4a2f4a3653349330a52c49b66fb52fb878b66fb5afb6efb1dda970b918b4afaeb92d49322536d437142a9231a5ab71252330252f4ab15db978bc3cbc3cb8d8b52fb2dd34d33754b46fb6afb3deb5efb25d30252c49b5afb5afb35db838b56f2d4931a5a1be38aa3c5532252e4a2c49384a3794384a3a4a33a6b938bb59bbd9b918b52fb42f302535132a92a1be1c8837943beb396ab05db66fb7b0aeb9b46fb1dda6e033a63a4a3d3631a531a5394a392a38ea37543ce53d153714b6afb978bbf9ba78b72fb35d252331a52a922e4a34d338ca39cab05db66fb35db72fb46f2a921c88388a3da63a8a3025396a384a382a379437d43cf53e963e563326b6afba58bc3cbad8b6efb4afb1ddaeb9a6e0b15db05d2e4a1c88b25dacb8b56fb66f2c4937943c753d3636933c153125b9f83453359336933c253c553e963ce52892b8b8bb79bc9cbbf9b8d8b72fb5afaeb9ab713326341330a5a1beafb9b3deab713513382a3beb3b4b3b0b3c45b52fba182a923613396a3dc6398a3ce53de63c552892b838ba98bc4cbc5cbad8b918b5efb72fb3de375439aa345338ea39ca39ca3754adb92e4a341332a6b0ddb6afb8583453398a3dc63e6638aa3aaa3d663e563c35acb8b5afb7f0baf8bc5cbb79b998bb59bc6cb8583593386a3b6b394a3225b35db938b5afb4afb4afb7f0b6efb878afb9;
    // label:6
//    input_ANN = 16384'h2a9237943d053c6537543653380a386a365335d338aa37943754390a3a4a39ea388a3a0a3c653cc53c453c353c553cc53c453c753cb53c353a0a3c953d053d05aeb938ca38ca3593341335d3365333a634d3359337943754386a382a394a3a4a392a3aca3c353cd53c653c353c653ca53d363d563c853b6b3a0a3c053c453c55afb93513ab712a9233a637d4365333a63593332635933693382a38aa38ea396a386a3a0a3c953d663cb53c253bab3b4b3c053b2b3b0b3b2b3b0b3bcb3c553c45ab71a6e0b15daeb931a537943453341334d32e4a3493345333a636d43794361338ca396a3cb53e163d563c953c353bab3a8a398a39ca3a0a3beb3c553b0b3acaa970a9702c49a1be332635932f4a2f4a302530252f4a2e4a31a5351337543653355337943a0a3d563d963c953c353cb53c353a8a3a0a3a0a3b2b3c053aca3a8ab15dadb935d3a1be2e4a33a62f4a2d492d492a922c492e4a31a533263754386a31a53326351339ea3c3539aa390a3b8b3b2b3b0b3aaa3a6a3a2a3a4a3a8a39cab62f30253693b05d28922d492e4a30a51c88a1bea9702f4a2a922c49341337543513345331a532253754380a37943aca3b4b3b0b3c053bcb3a8a3a2a3a0a396ab4ef38ea30251c882c492c492f4aa1beadb9a1beacb8252328922f4a302534d334d3332630a53225341339aa386a3a6a3beb3bab3cb53c453aeb3aaa3a0a39ca30a534132f4a31a52c492e4a2c492892adb9a6e02e4a2e4a2892332634d3365336933794351334132f4a369330a5388a3bcb3c153b4b3a6a3a8a3a2a3a2a39ca302532a635532c49a1be1c88a1be31a52c49a970aeb9a9702c493225349331253453388a38aa351331253513289236133c253bcb3a8a3a4a3a8a39ea3aaa39ca36d43aca31a5a9702892acb8a6e0ab71adb9afb9adb925232f4a2e4a2a92b4efadb93653394a37d435d335d3341338aa3d263beb3bcb3c153b8b3a8a3a0a39aa3dd63ca5a970349337542523b0ddb05dafb92f4a2d49b15db838b52f31a5adb9b2dd33a638ca36133613371438ca3cf53d763c153bcb3c053bcb3b0b3a8a39ea3e163c05b46fa6e0b3deb770b3deafb9ab7134532c49b66fb9d8b46f30a5398a3beb388a396a3693332637d43a0a3ce53d863d153c753c453c253b0b3aeb3aaa3e963b0b28922523b7b0b62fb46fb3de2e4a3513b35db7f0b5afa6e0a6e02f4a3a4a322532a634d32c49388a3b6b3d263de63d763cc53c653c253bab3beb3b6b3b0b398a3a4a3225b66fb4efb0ddb46facb8adb9b838b72f1c883125b05db62fb42fb7b0b42fb5afa1be382a3a8a3d153d263d263c753b2b3c153c053c553c15384a3b2b3c053225b6efb66fb0dd1c88b3deb6afb8d8b8d8b818b15db4efb858b838b72fb770b7f0b05d2f4a398a3c853cf53d763beb3794398a3c753c753c353794392a3b0b3553b4efb42facb83453b0ddb898b9f8b7b0b878b2ddb25db838b6efb56fb52fb66fb6efaeb93aeb3d153e463df63a8a359333263c253d363c453794375437d42e4ab4afb5afb52f35532892ba38adb93453b56fb46fa1be2a921c88b15d1c882a9231a5390a3d763ea63f063e563aca35d330253a0a3da63cf535d33613392a2d49b770b6afb4ef371438cab93831252892b918b05d39ca36d439ea365338ea3beb3ca53e463ed63e563e963d863b2b3025252337543dd63d863513382a3b4b32a6b72fb858b72f31a53db62c49b5afb2ddb62f30a5382ab8381c88390a3beb3da63dc63e763da63cf53e163d263aeb2e4ab5af2f4a3df63e26349335d337543025b5afb818b62f30a53f563e56375432253125384a396aafb9b4af36933ca53e263cf53ce53cc53ca53e563e063b4b1c88b818b4af3cb53e2630a5322537943553b3deb56fa6e038ea3f263f763ec63de63cb53c253cd53aaa386a3a2a3c653e563e263e063de63cb53d463d263beb32a6b6efb6af3b4b3e262c49322538aa37141c88b05d32253b6b3d053bcb3d863ea63e763d863cd53a8a3c853e263dd63e863ec63ee63f463e263cd53ca53c2539cab05db46f398a3e062f4a3714369335133413a1be3225379436d43a8a3c353bab3b2b3b8b39ca3beb3e863fc63fd63f863f463f163fc63fa63eb63df63c353c153754b0dd36133db6369339ca34d32a92361335d3b0ddb5af2d493bcb3a0a3a0a390a39aa3aca3c453d763eb63f063f663f763fb63fb63f663f963db63beb3d563c7535132d493aeb365335d3341334533553388a34d3b05db3de34d31c8836133a4a396a38ea3a0a3bcb3d263da63e763ee63f663fb63f263f063d863d153eb63d863c6538ea36533653359334d334932c4930a537d43a0aadb9349339ca394a3a4a35d33453386a3a2a3bcb3c653cd53cc53d663e163d663d363d963db63d663bab388a3ce53b4b3754355338ca384a2a9230a535933a2a37d431253aca3a4a39aa35d3349336933a4a3a6a39ca3a0a3b0b3beb3bcb3a0a3a6a3b8b3bab3b4b39ea37943c753c15351335533a8a392a31a536d4390a38ca382a3a4a398a34d337943653355335d338ca388a384a39ea3a6a39ca392a37d4388a38ca392a394a3aca3c553aaa3693396a382a388a33a63493361336d4365332a637d436d4341336933613361336533754384a398a3b0b396a386a382a3693361337d437d4386a3aaa3aaa382a34d3382a351330a5289234d33513349334d333a6332630a5312535d336d438ea39aa388a390a392a398a392a380a37943653345336d43714386a394a396a380a36d4361330252a9232a638aa3a8a38ca3613355338ea375436d4371436d4398a3b6b3a0a390a380a388a386a3653369335533413361337d436933653375436d43794;
    // label:1(��ȷ��)
//    input_ANN = 16384'h3c053a4a38aa386a369333a632a633263125332635d3379437d4375437d432a63a2a355338ca2c493a8a3b0b3c253c653d963d153c953d763d863dd63df63df636d4351334133693369334533513a9703613371438aa396a39aa394a394a3a8a3b4b3b6b3bcb3c753c453c853d053ca53cc53ce53e863e563d863da63dd63de63453351335132c49388a37d4386a32a6396a39ca3a6a3b0b3b6b3aeb3b0b3bcb3c353c553c853cf53cc53c953ce53d053cc53e363fd63f263db63d863dc63dd6380a388a380a386a382a39ca3a4a3b0b3b4b3b6b3bcb3c253c453c153c353c653ca53cb53cc53cc53ce53d053ce53cf53d963ef63f763ec63d763d763dc63dc638ca392a37d438aa39aa3b6b3bcb3c353c553c653c853cb53cb53c953ca53ca53cd53cd53ce53cd53cf53c253a2a3cf53e563e863ef63dc63d363cf53d863db6396a39ca3aca3c253c953c853c853cc53ce53ce53cd53ce53ce53ce53cd53cb53cc53ca53ca53cb53c75379438ea3c853d563e363df63c753c553c353d663da63c853cd53d053d263d153d153cf53d263d153d153ce53cc53cd53cb53ca53c653c853c853c853ca53b4b392a3d263e363cb53d663ca53c353c853cc53d863d863d963d763d763d563d053d153cf53d263cf53cf53cb53ca53ca53c653c653c053c253bcb3b4b3b8b3aaa3c753f663fa63d863cb53cd53ce53d363d363d863d863da63d663d463d463d053d153cd53cf53cd53cc53c853c653c353a8a3a8a39aa3a2a3a2a3a8a3aeb3b6b3dd63f763f463d663cd53cf53d053d363d463d763d963d763d563d363d363cf53d153cd53cd53cd53cb53c453aaa39ea38ea3a2a3a4a3b0b3bab3b4b3aca3c253d363d763d863ca53cb53d363d153d563d563d763d963d563d463d153d263cf53d153ce53ce53cd53cb53c253aca3beb3a2a3a4a38ea3326b35db978bb393125384a3bab3e363c753c153d053d463d663d663d963db63d263d263cf53d153cd53cf53ce53ce53ce53c953c953beb384ab62fba38bb39bc6cbc5cbc4cbb99b8b8bc3cb3de3ea63ef63e163aeb3c953d963d963db63dd63d053d153ce53d053cc53cd53ce53cd53cf53ca539ca3025b42fb56facb83493380a39aa3bab3c9534d3bdddbcac3a6a3f963fe63d153a6a3d763db63dd63df63cf53d053cc53cf53cc53cc53d053ce53cf5394a355338ca3a4a39ca3d363f463f263e063f563f6631a5bd3cbd5db56f3e2640033f263c953da63e163de63e063cc53ce53c953ce53cc53cc53d663d263b2b38ca3c553d563c253aeb3d663ef63f963da63e963c05ba78bcdcbcacbc7c37d43f763f663f063e963e763e263e163cb53cf53c953cd53cd53c653a8a3b6b39ca3cf53ca53c4539ea3b4b3da63e263e463beb3326bb18bd2cbcccbd0cbc7c34d33cc53ed63f863ea63bab3bcb3e363cc53d053ca53cd53c953c053754384a3b6b396a3ca53c553aaa3c1539eab62fbb79bd6dbebdbebdbd9dbd9dbd4c34133de63c053ea63fa63c15adb930a53e163cc53cf53cc53cc53c953d463d053c253a0a3aca3e563e263da63e96b15dbf1dbebdbe9dbe0dbd9dbd9dbdadafb93df63ed63da63d153c052523b6efb56f3d463cd53d053d053c5537143c053d863d053bab3e263ef63ed63d153d86b6afbd9dbcbcbc2cbc1cbd0cbdbdbdcdb8183a6a3c25388a2a92b3deb46fb3deb6ef3c853d053d363c75adb9b9983a0a3e263db63c953f063fa63f163c853b6bb818bc6cbb99bb39bc8cbcccbc3cbcfcbdbdb978b46fb7b0b6efb62fb4afb35da6e03d663d153d963493bd9dbab837543d963d963cf53fc63fd63fa63ea63c95b8d8bc0cbad8bbf9bb9932253b4b388ab858bc8cbbb9b9d8b8d8b7b0b4afacb83b8b3f063d663d26aeb9b7b0b25d32253d153d463e9640233fd63f363dd63c35b918bb59ba58bc2c33263ee63ee63eb63d05b62fbc0cb9d8b4efb05d1c883c353f763f063db63c7539aa3e663aca31253ca53d263f4640033f863c2537d43593b978bad8baf8b9983d863e863d663dd63f463b4bb5efb1dd2e4a30253c753fb63fb63e863dc63cb53ca53e463c352c493b4b3e363f963f763e763a4a394a32a6bc1cbc1cbc5cb2dd3e863db63e763e963e863e8634d3afb91c8838ca3f063f863e963df63e063da63cb53c553c252d493a2a3e663f363e263cb53a6a3a8ab35dbc3cbb39bb5930a53e363cf53d053db63eb63f863b4bb0dda1be3c553f763ef63e563e063e863e463d363c853c4532a63a6a3ec63ec63ce539aa36d43693b5efb958b938ba1831a53e063cb53b8b3d263e263f763db6341336d43e163fe63f663f063e963e963e563d763ca53c3535d3384a3cd53b6b34d3b4afb998b9d8baf8bbb9bb99bb7925233de63cb5384a38aa3d263eb63f363b4b3c453f86401b3fc63f663ec63e463e363dd63beb3beb386a3aca3ce53c653b6b39ea38ca382a369336533714371439ca3e263c653c753c553e763f0640033f363fa6401340033ff63fa63ec63e163da63dc63dc63da63dc63f3640033ff63ff63fd63fc63fb63f863f763f763f863f863fe63c453c253d663ce53f76402340234023401b400b3fe63f963ec63d863d263d363e263f063f763f063e963f263f563f263f263f263f463f563f863fc63fd640033ef63c853bcb3dd63ff640234013401340133ff63fa63f063e963d863d563d463d263ce53c953b6b3bcb3df63e763df63dc63da63de63e363e663eb63ee63f363f863f063ee63fd63ff63fd63ff63fe63fd63fa63f563e963e963d563d363c653a2a37943794390a3b6b3d563ce53c853c753c453c453c653c853cf53d763df63e163db63dd63f063f763f563f363f363f663f263eb63e763ea6;
    // label:6
//    input_ANN = 16384'h39aa39ca39ea3a6a3a2a39ea392a390a390a38aa37d4390a39aa3a4a3a8a3aeb3bab3c053c253c353c653c953cd53d263d763dc63e063e263e163e763ec63f06398a39aa39aa3a6a3a4a3a2a394a38ea394a398a388a386a39aa3a4a3aca3b0b3b6b3beb3c353c153c653cd53cf53d563d963de63e163e363e263e863e963e8639ca39ea3a0a3aaa3aeb3a0a398a3b2b3a4a39ca398a382a37d4398a3aeb3b0b3b6b3c053c553c453cb53cf53d363d963db63de63df63dc63d863d963d763d5639aa39ea3a0a3a4a3b0b39aa3a8a3d2639ea386a39aa392a37143794398a3aaa3bcb3c753c753c753cc53d053d053cf53cc53ca53c653c453c353c553c753c853a0a3a2a3a2a3a2a3b0b3a2a3b0b3cd53a2a3a0a3b2b3b4b3aca396a394a39ca3a8a3c553c453c153b4b3b6b3b0b3aaa3aaa3aca3aaa3aaa3aca3b4b3beb3c653a8a3aca3aaa3a6a3b2b3b6b3bcb3bcb3bcb3bcb3bab3b6b3b2b3aca3aeb3aaa39ca39ea390a38ca38aa388a38ea38aa394a39ea39ca3a4a3b2b3c053c753ce53aeb3b0b3b4b3b0b3b2b3ca53de63d463bcb3bcb3bab3b6b3b2b3bab3aeb39aa39ca394a371435d3382a388a384a382a396a3aaa3b0b3b8b3c253c653cb53ce53b4b3b2b3b4b3b0b3bcb3d053e163df63c753c453c453c353c453c053aeb39aa390a3a0a39ca384a37d436d43714398a3a8a3aca3b0b3b8b3beb3c153c453c853b4b3b2b3aeb3a0a398a382a3a6a3da63c953c453b4b3a0a3a4a39ea39aa3a8a398a394a39aa39ea38ca382a379438aa3a2a39ea3a4a3aeb3b4b3bab3b8b3b4b39ca38aa35d33125ab71b4af382a3d663c753c253aeb382a379435d3379439ca398a392a392a398a396a38aa3794369338ea396a39aa39ca39aa39aa39aa39ea2f4aacb8b3deb5afb6efb7b03a2a3d663c153c753cc5394a371434533553394a394a390a396a394a394a396a38ea382a388a388a37d4382a386a38ca390a398ab42fb56fb62fb6afb6efb72f398a3dc63bab3b8b3c75398a365338aa3714388a396a38ca392a398a390a394a39ca38ea392a38ca37143754380a386a38ea39aab4efb5afb62fb56fb4efb4af35133d963c35396a38ca36d432a63794388a384a394a380a38aa398a392a38ea3a2a39aa382a390a382a36d43794388a39aa3acab35db35db2ddb15db0ddb05d25233b6b3dc63c1538ea371434133413386a388a390a3714384a390a390a390a3a0a3a4a3754388a390a380a38ca39ea3b4b3c45ab71ab71acb8acb8aeb9b15db25d2c493a4a3c553d663c8539aa38ea396a38ca382a36133613380a38ca390a3a0a3a6a38ea384a3a4a398a3a2a3bab3c553c65a1bea6e0acb8afb9b3deb5afb3deb15db3de36133d563d05386a38ca396a386a3613322533a63553382a392a39ca3a0a3a2a386a3aaa3b6b3bab3bab3b4b3acaab71b15db42fb5afb6afb5ef252335d3b46facb83326380a34d3351338ca388a3714349334533593380a392a396a398a3a8a38ea39ea3aca39aa39ea3a4a3babb35db4afb56fb62fb7b0b918b8d830a5b8f8bb79b2ddaeb937d4a1be3413388a37143613351335d337d4386a38ea392a3a6a398a390a39ea392a3aca3cb53d96b4efb6efb8f8bb39bd2cbe4dbeedbb99b56fbc0cb858b918386a25232e4a380a379436533593359336533714382a38ea39ea39ea390a3b6b3c453d153d963d86baf8bcccbe0dbeedbf3dbebdbf1dbecdb6efb6afb838bad836d4369328923693380a36533613361335d335d33653388a398a3a2a3a2a3ca53d563d663d763d56beddbf3dbf3dbf4dbe9dba38ba78bc4cb42f1c88b35db4af3493375430a535d3371435d335d33593355335533653388a39ca3a8a3aeb3c353d263d263d463d66bf3dbf3dbf3dbf6dbe1d3025365333a6355331a5332635933714379437d4388a36d43553355335933553369338aa396a3a6a3b2b3b0b3a6a3c353cf53d153d46bf2dbf2dbf0dbe5dbc1c312534933225386a390a39ca3a0a39ca396a3b8b3c75392a37d43794382a388a38ca386a384a396a3aaa3b8b39ca3a0a3cb53d153d15be9dbd3cba78b52fadb9a1be25232523380a3c553c553c153b8b396a390a3d053d463bab3aeb3a0a38ca3794369337d439ca3bab3bcb3a4a390a3bcb3d053d05b62fa1be2e4a3025302532a63613380a379439aa3c753cc53bcb382a37943aca3c653b2b3a0a394a37543613365335d3384a3c053c153bab39ea398a3c353d05359334d334533593380a38ea386a379435d33513380a3a6a39ea38aa390a39ca3b6b3aaa394a388a33262e4a34d33693369338ea3beb3c053b8b394a3a4a3cf53754388a392a396a388a379436d43714380a392a3a0a3a8a3c453c253a4a392a3a6a3aca398a388a3125252334533794386a38aa3a8a3bcb3c153aca39aa3c353a2a3a4a396a38aa37943754386a39ea3b6b3c753c253a0a3b4b3c853bcb39ea3a8a3b2b3a8a3a8a390a3653375438aa392a394a3b0b3c453c353c153b0b3aeb39aa394a38ca38ea398a3a6a3c053ca53ce53cd53bcb39ca3a6a3bcb3a6a3bab3c553c753c553c553c653b0b39ca392a396a3a8a3c653cb53c753c753c653b8b390a398a3a8a3c053c853cb53cd53d053d053d053beb3a0a3a6a3aeb3b0b3c853c953ce53ce53ca53cb53c953c153bab3bcb3c453ce53d053cc53cb53cf53cb53b8b3c753d153d663d363ce53ca53cf53d053d363c453aeb3aeb3a8a3c453c953ca53d053cb53c853cd53d153cd53d053cf53cc53d053d363d263d053d363d663d963dc63d863d963d263d263d363d263d153d563c753b0b3bcb3aaa3c553cf53d053d263d053cd53cf53d263ce53d153d263cf53d263d663d963d663d663d96;
    // label:8����ȷ�ģ�
//    input_ANN = 16384'hba18b9d8b66fb46fba98bc3cbc7cbcccbd0cbd3cbd5dbd0cbdbdbdedbe1dbe4dbd3cbe0dbe5dbe7dbe8dbe5dbe7dbe7dbe9dbdedbe2dbeadbe4dbdedbe7dbe9dbb59bb59b878b52fbb59bcccbcecbcfcbd4cbdbdbdbdbd2cbe0dbe5dbe6dbeadbd8dbe1dbe5dbeddbefdbe4dbe6dbecdbecdbe0dbe6dbefdbe4dbe0dbeedbefdbb99bb79b8f8b5afbbb9bd0cbd4cbcbcbd3cbdfdbd9dbd2cbdcdbe1dbe1dbebdbd9dbe0dbe5dbeadbe2dbcecbe2dbe9dbefdbe1dbe8dbf2dbe6dbdedbf2dbeddbbd9bb79b8f8b66fbbd9bcecbd6dbcfcbd5dbe1dbdadbd1cbd5dbe0dbdadbebdbdbdbdedbe4dbe1db9d8b8d8bdddbeadbf0dbe0dbe6dbf2dbe5dbdbdbf0dbebdbc3cbc0cb958b5afbbd9bcccbd7dbcccbcecbe3dbd9dbcfcbd2cbdedbcccbe4dbdbdbd9dbe3dbd5db7f0b8b8bd9dbe5dbefdbdfdbe3dbeedbdfdbe0dbeedbe8dbc5cbc1cb998b42fbbf9bc9cbd8dbcecbd1cbe4dbd6dbcfcbcfcbdcdbbf9bc5cbc8cbc7cbe6dbc1c3326b770bdadbe0dbeddbdddbd9dbe7dbdadbdedbeadbe1dbc3cbbb9b958a970bb39bc2cbd5dbcecbd3cbe0dbd0cbcccbcfcbdcdba98b918bab8bad8bcacbaf83025b1ddb998ba98bd6dbd7dbcecbdedbd4cbd7dbe4dbdadbc5cbbd9b8f8acb8bb99bc8cbcbcbcacbd2cbdadbcacbcccbcecbd0cbbf9bc5cb918b15d3653398a3a8a3b6b3b6b3c453714b9f8bc6cbd7dbcacbc0cbd9dbd1cb8d8b838b52f1c88b838b938b770ba18bb79bbd9bb39bbf9bc2cbb39bb18bb99b35d345337d43794384a386a37143b4b3aca32a6b62fb938b770b42fbb39b97834d334933513379436d4365335d33025a1beab71afb9b2ddb46fb0ddb52fb5af2c4934d334d334d337d437d4388a398aaeb92f4ab42fb1dd35d337142d4933263b6b3a4a3a6a3b2b390a382a392a38aa388a369337543693359334932e4a3225379437943754382a398a3a8a375434132c493613b05dbb1833263693386a382a3c253aca398a394a3125341338ea3b0b382a30a53693365330251c882e4a345334d3361335d335933714388ab52fbab8b9b8b1dd3693bbd9b2dd384a38ea38ea3b6b380a369339ca359335d339aa388a2523b25db0dd30a531252a9233a636d4382a382a36d43493359331a5b8d8bb59bc6cbad833a6b72fb8383aeb390a390a394a3754380a39ca390a3aca3a2a38ea375433a61c882d4932a6302530a534133453332633a62d492d49b3deb9b8b9b8ba58ba38b46f3125b6ef3b2b3c253a8a38ca38aa388a394a394a3a2a3a2a37d43025ab71b1ddb46fb5afb5efb56fb42fb7b0b818b770b770b5efb818b938b8f8b958b858b7b0388a39ea3c053ca53c053453355331a533a631a5b15db35db56fb72fb898b8f8b8f8b958b958b998b838b838b8d8b898b56f30a52a92afb9b6efb878b72fb7f036d43c1538ea39ea3b0b2e4a32a62523b25db0ddb42fb6efb72fb7f0b878b8f8b938b978b958b8d8b770b1ddb2ddb3dea1be386a3413b05db52fb7b0b6efb6ef1c88b0ddba98b46f371434132d49a970302535933613b2ddb7b0b878b898b898b818b62fb42fb15db05dab71b15db770b56fa970b3deb72fb5afb6afb4efb52fb3deb5afb5efb46fb1dd31253653394a39ca37542c49b05db62fb770b46fb05dacb8aeb9b1ddb46fb5efb770b52fb72fb838b5efb6efb818b72fb5efb56fb56fb15d2a9233263125b35d36d43aca396a2c49b3deb66fb42fafb9a9702523afb9b4afb6afb838b878b7f0b6efb3deb5afb770b66fb62fb6efb7f0b56fb2dd2e4a365338ca3aeb398aa6e02f4a30252d49a970a970a970b0dda9702523b52fb6efb770b6efb62fb25d2c4935d3380ab05db66fb66fb66fb5afb3de31253794388a39ea3bcb3b4b3b0b3c0530a52523a970a6e0a970aeb9b15db15d1c88afb9b05db2ddb42fb35d37543b8b3c053c152f4ab62fb35dacb831a5375438aa390a3a4a3c053c053aca3cf53e7639ea2d49aeb9acb8acb8acb831a53613382a38aa390a2d49b42fb2dd361339aa38ca386a332633a63693384a38ca38ea3a8a3bab3c753cd53c853d363e363e963aeb34132e4a2f4a2c4930253a0a3beb3b2b3a6a3a0a3025b35db1dd2e4a35d3382a394a396a394a392a38ea39ea3beb3cf53ca53cf53d263db63e363e663e963a4a361331a530a52c492a92386a396a37d43653341332a63613392a3aca3b0b3a4a39ea392a38ea3a0a3c353cb53c953c053c753d663db63de63e363e663e863a0a37143125322533a634d3375438aa394a3a4a3b8b3beb3c053b6b3aeb3a2a39ca3a6a3b4b3c353cb53cb53c953ce53c553cf53df63e163e063e363e663e363beb3b8b3aaa3bab3c153c653cb53cc53ca53c653c253beb3b6b3b2b3b4b3bab3c453d153d463c853c953cb53d363d863d463dd63e263e163e163e363e263e363dd63df63e263e063da63d863d763d263c853c553c453c653cb53d153d263d153d463cd53aca3c253d263d763da63da63de63e263e363e263e163e063df63eb63de63e163e563e363df63dc63db63da63d763d863db63db63d763d153ce53ce53d363c6539ca3c953de63db63d963e063e263e363e263e063e063db63e863f663e163e263e663e563e463e263e263e063de63d963d463d263cf53cf53d053d363db63cf53aeb3d563e263db63e363e463e463e463e263e063de63df63fb6400b3e863e463e663e263df63dc63da63d763d563d363d153d363d363d563d963de63e863da63bcb3d863e063e363e463e463e563e563e663e163dc63f364013400b3e163df63dd63db63db63da63da63d963d863d763d963dd63e163e763f063f763ff63ee63cc53dd63e763e663e663e563e663e863e863dd63e96400b401b3ff6;
    // label:3
//    input_ANN = 16384'h3f263f263f563d36ab71b52fb46fb35dafb9b05db42fb3deb35db2ddb2ddb3deb25d2523380a3b4b38ca38ca1c88b858b6efb7b0b72fb7b0b7f0b770b6efb66f3f263f363f463e462e4ab858b6afb46fb05dacb8b0ddb52fb5efb56fb46fb52fb6afb4ef32a63b6b3c45394ab66fb9b8b918b978b958b978b958b8f8b898b8783f263f263f263ef636d4b858b56fb15db15db3deab71afb9b5afb5afb56fb6afb818b8f8b7b035933c95384ab9b8ba98ba58ba58ba18ba18b9f8b998b938b8d83f263f263f163f463a6ab62fb1dda6e0b56fb770b5afa6e0b52fb858b8b8b978b978b998b81831a53a2aa1bebbd9bbd9bb39bab8ba58ba58ba78ba58b9d8b9b83f063f263f163f363cb5b05da6e03025b6afb998b9b8b25d1c88afb9b46fb878b978b8f8b5af31253613b7f0bc5cbc9cbc9cbc3cbbd9bb99baf8ba98ba18b9783ef63ef63ef63f063de633a6a1be2f4ab46fbab8bbb9b66f332635d335d3a1beb35db25d25232523afb9b9b8ba78bb99bc5cbc8cbc4cbc9cbc9cbc3cbc1cbb993ed63f263f063f163e763553b6efb42fb52fbad8bbb9b8b82c49382a3693349336d433a636132c49b978bc1cbab8bb99bc7cbc9cbc9cbcfcbcfcbcdcbcecbd1c39ca3dd63ee63e8638eab898ba38b52fb42fba38bb18bab8b7f0a1be2a9232a638ea361335d32f4ab9f8bc5cba38bc6cbe1dbdbdbe1dbdcdbc4cbc9cbd2cbd9db8f8b42f36d434d3b8b8ba78b9d8b25d3225b770baf8bb59ba78b918b56f1c883413341332252c49b838bbb9ba38bcfcbe2dbdbdbdadbc9cba38bb79bd5dbdedbaf8ba58b8b8b998bab8baf8bab8b0dd3453b52fb998ba38ba58ba58b818aeb93794332632a630a5b6efbab8bc5cbdedbdfdbe2dbdfdbbd9b9d8ba18bc5cbe0dbbb9bad8b9b8ba58bb99bc2cbab8ab71a970b818b978b9f8ba58b958b5af302536533326332632a6b62fb918bc2cbe4dbe9dbe9dbe5dbc5cba38ba38bb18bd3cbbf9bbf9baf8ba58bbf9bc5cba58b1ddb56fba18ba78ba38ba58b6efa1be36533453a1be30252e4ab66fb878ba78bdfdbebdbe9dbe4dbcfcba58ba18ba38bb79bc0cbbd9bb59ba78bb39bb59b9d8b7f0b66fb898b958b7f0b7f0b770aeb93225a1beb66fa6e0b25db72fb7f0ba78bdcdbe8dbebdbe9dbdcdbc0cba58ba38bb18bc4cbbb9bb18b9f8bb18b7f0b5efba98b6afb1dda6e0a6e0b6efb66facb8b1ddb818b770b2ddb6afb4afb56fbb39bdadbe7dbeadbecdbe9dbdadbb18bbb9bcfcbc6cbbf9bb59b9d8bb39b25d2523bbd9b9d8b978b818b818ba58b8982a923413b858b858b35db5afb898b8b8ba98bdddbe7dbe8dbe9dbf0dbe6dbc2cbcecbdbdbc7cbb59bb39ba18bb39b4af31a5bbd9bc0cbaf8bad8b9b8b7b0b838b6afaeb9b3deb938b66fb15dba38b938b818bb79bdedbe6dbeadbeddbd7dbcfcbdddbdcdbcbcbb39b938b8b8b9b8b7f03225b998bc9cba78b838b978b838b56fb838b8183513b46fb978a1beb56fb898b15d3794b15dbc8cbe3dbe1dbc5cbcfcbe4dbdedbcdcbbf9b72fb52fb7b0b938b66fb838bc3cbc6cbc1cbcacbab8b858b898b77034d33225b918ab71b35dbab8b5af3453384a2892b938ba58b9d8bc7cbe5dbe1dbcfcbc7cb8b8b5efb918ba78ba98b9b8ba98bc7cbcdcbd6dbd5dbbf9ba58b8b8aeb93714b46fb05db4afb998b46fb42fa1be34d3acb8b56fb3deb918bcfcbdfdbd1cbcacbb18b8f8bb39bb79bb79bc2cba18ba18bb18bc0cbc5cbc9cbc2cb958b898a9702c49b6afb878b5efa1beb2ddafb92c49b46fb6efb35db15db5efbb99bd3cbcecbc2cb998bab8bbf9bb18bb79bbb9ba98bad8ba78b898bb59bc0cbb39bc8cbb59b42fb8b8b72fab712f4ab1ddb25db4afb770b56facb8acb8b05db4efbd1cbcfcbc9cba38b938bb79bc1cbaf8bc0cbc6cbc7cb978b46fb958ba38ba18bbd9bbd9b938b838a9703025adb9b3deb56fb770b5afafb91c88afb9afb92f4abcecbcdcbcecbb39b7f0bb18bcbcbc9cbc5cbc8cbc7cb9f8b5efb8d8b9f8b998ba18b9f8b978b4af35132f4ab46fb52fb52fb770b5afaeb9aeb92a9234133653bcdcbc9cbcbcbc2cb7b0ba98bcbcbcfcbcfcbcdcbc1cba98b978ba78bab8ba38bab8ba38b8f8a6e03453acb8b56fb46fb42fb8f8b6efb35db25d3025341332a6bcbcbc6cbc6cbc2cb8d8ba78bc7cbc7cbc7cbc7cb9f8b25db8d8bbb9bab8ba58ba98ba18b6af25232e4ab05db46fafb9b0ddb7f0b66fb46fa6e01c8825232f4abcacbc4cbc1cbb39b9b8ba58bc5cbc5cbbf9bbd9ab71394ab4afbb99ba58b958b958b838b3de1c8831a5aeb9b15dab71adb9b15db05dacb8a6e0a6e0312534d3bcacbc2cbbd9ba78b8d8b938bc3cbcacbc4cbb79acb838cab46fbab8b8d8b770b770b46fadb931a53413ab71acb82d49a6e0302534d330a5aeb9acb81c882a92bc9cbbf9bb39b9b8b818b818bb79bcccbc8cbb18b818b4efb978b878b5afb4afb15da9702c4937d4349325232c4930252d49345335d334532523b25db25dadb9bc6cbaf8ba78b938b66fb5efbad8bcacbc8cbb18ba18ba18b8f8b56fb0ddb0ddab712d493513390a32252d492d492c492d493453369333a6a6e0b25db0dd2892bb18b8d8b8d8b978b5afb05db978bc4cbc5cbb59ba78b998b838b35da970aeb92c49341338ca386a3225341331a52a922a92349334932d49a1be1c8825233025b898b52fb72fb958b7b02892b4efbb99bc1cbb59bb18ba18b25d34933593332632253653394a35933493351331a51c88302530a52c492f4a332630a52523a970b3de2523b05db4efb5af31a53025b958bb18ba18b918b52f35133a0a3b6b39ea37d438aa37d435933653361331252e4a312530a53513361334531c88adb9a1be;
    
    
   input_ANN = 16384'hba18b9d8b66fb46fba98bc3cbc7cbcccbd0cbd3cbd5dbd0cbdbdbdedbe1dbe4dbd3cbe0dbe5dbe7dbe8dbe5dbe7dbe7dbe9dbdedbe2dbeadbe4dbdedbe7dbe9dbb59bb59b878b52fbb59bcccbcecbcfcbd4cbdbdbdbdbd2cbe0dbe5dbe6dbeadbd8dbe1dbe5dbeddbefdbe4dbe6dbecdbecdbe0dbe6dbefdbe4dbe0dbeedbefdbb99bb79b8f8b5afbbb9bd0cbd4cbcbcbd3cbdfdbd9dbd2cbdcdbe1dbe1dbebdbd9dbe0dbe5dbeadbe2dbcecbe2dbe9dbefdbe1dbe8dbf2dbe6dbdedbf2dbeddbbd9bb79b8f8b66fbbd9bcecbd6dbcfcbd5dbe1dbdadbd1cbd5dbe0dbdadbebdbdbdbdedbe4dbe1db9d8b8d8bdddbeadbf0dbe0dbe6dbf2dbe5dbdbdbf0dbebdbc3cbc0cb958b5afbbd9bcccbd7dbcccbcecbe3dbd9dbcfcbd2cbdedbcccbe4dbdbdbd9dbe3dbd5db7f0b8b8bd9dbe5dbefdbdfdbe3dbeedbdfdbe0dbeedbe8dbc5cbc1cb998b42fbbf9bc9cbd8dbcecbd1cbe4dbd6dbcfcbcfcbdcdbbf9bc5cbc8cbc7cbe6dbc1c3326b770bdadbe0dbeddbdddbd9dbe7dbdadbdedbeadbe1dbc3cbbb9b958a970bb39bc2cbd5dbcecbd3cbe0dbd0cbcccbcfcbdcdba98b918bab8bad8bcacbaf83025b1ddb998ba98bd6dbd7dbcecbdedbd4cbd7dbe4dbdadbc5cbbd9b8f8acb8bb99bc8cbcbcbcacbd2cbdadbcacbcccbcecbd0cbbf9bc5cb918b15d3653398a3a8a3b6b3b6b3c453714b9f8bc6cbd7dbcacbc0cbd9dbd1cb8d8b838b52f1c88b838b938b770ba18bb79bbd9bb39bbf9bc2cbb39bb18bb99b35d345337d43794384a386a37143b4b3aca32a6b62fb938b770b42fbb39b97834d334933513379436d4365335d33025a1beab71afb9b2ddb46fb0ddb52fb5af2c4934d334d334d337d437d4388a398aaeb92f4ab42fb1dd35d337142d4933263b6b3a4a3a6a3b2b390a382a392a38aa388a369337543693359334932e4a3225379437943754382a398a3a8a375434132c493613b05dbb1833263693386a382a3c253aca398a394a3125341338ea3b0b382a30a53693365330251c882e4a345334d3361335d335933714388ab52fbab8b9b8b1dd3693bbd9b2dd384a38ea38ea3b6b380a369339ca359335d339aa388a2523b25db0dd30a531252a9233a636d4382a382a36d43493359331a5b8d8bb59bc6cbad833a6b72fb8383aeb390a390a394a3754380a39ca390a3aca3a2a38ea375433a61c882d4932a6302530a534133453332633a62d492d49b3deb9b8b9b8ba58ba38b46f3125b6ef3b2b3c253a8a38ca38aa388a394a394a3a2a3a2a37d43025ab71b1ddb46fb5afb5efb56fb42fb7b0b818b770b770b5efb818b938b8f8b958b858b7b0388a39ea3c053ca53c053453355331a533a631a5b15db35db56fb72fb898b8f8b8f8b958b958b998b838b838b8d8b898b56f30a52a92afb9b6efb878b72fb7f036d43c1538ea39ea3b0b2e4a32a62523b25db0ddb42fb6efb72fb7f0b878b8f8b938b978b958b8d8b770b1ddb2ddb3dea1be386a3413b05db52fb7b0b6efb6ef1c88b0ddba98b46f371434132d49a970302535933613b2ddb7b0b878b898b898b818b62fb42fb15db05dab71b15db770b56fa970b3deb72fb5afb6afb4efb52fb3deb5afb5efb46fb1dd31253653394a39ca37542c49b05db62fb770b46fb05dacb8aeb9b1ddb46fb5efb770b52fb72fb838b5efb6efb818b72fb5efb56fb56fb15d2a9233263125b35d36d43aca396a2c49b3deb66fb42fafb9a9702523afb9b4afb6afb838b878b7f0b6efb3deb5afb770b66fb62fb6efb7f0b56fb2dd2e4a365338ca3aeb398aa6e02f4a30252d49a970a970a970b0dda9702523b52fb6efb770b6efb62fb25d2c4935d3380ab05db66fb66fb66fb5afb3de31253794388a39ea3bcb3b4b3b0b3c0530a52523a970a6e0a970aeb9b15db15d1c88afb9b05db2ddb42fb35d37543b8b3c053c152f4ab62fb35dacb831a5375438aa390a3a4a3c053c053aca3cf53e7639ea2d49aeb9acb8acb8acb831a53613382a38aa390a2d49b42fb2dd361339aa38ca386a332633a63693384a38ca38ea3a8a3bab3c753cd53c853d363e363e963aeb34132e4a2f4a2c4930253a0a3beb3b2b3a6a3a0a3025b35db1dd2e4a35d3382a394a396a394a392a38ea39ea3beb3cf53ca53cf53d263db63e363e663e963a4a361331a530a52c492a92386a396a37d43653341332a63613392a3aca3b0b3a4a39ea392a38ea3a0a3c353cb53c953c053c753d663db63de63e363e663e863a0a37143125322533a634d3375438aa394a3a4a3b8b3beb3c053b6b3aeb3a2a39ca3a6a3b4b3c353cb53cb53c953ce53c553cf53df63e163e063e363e663e363beb3b8b3aaa3bab3c153c653cb53cc53ca53c653c253beb3b6b3b2b3b4b3bab3c453d153d463c853c953cb53d363d863d463dd63e263e163e163e363e263e363dd63df63e263e063da63d863d763d263c853c553c453c653cb53d153d263d153d463cd53aca3c253d263d763da63da63de63e263e363e263e163e063df63eb63de63e163e563e363df63dc63db63da63d763d863db63db63d763d153ce53ce53d363c6539ca3c953de63db63d963e063e263e363e263e063e063db63e863f663e163e263e663e563e463e263e263e063de63d963d463d263cf53cf53d053d363db63cf53aeb3d563e263db63e363e463e463e463e263e063de63df63fb6400b3e863e463e663e263df63dc63da63d763d563d363d153d363d363d563d963de63e863da63bcb3d863e063e363e463e463e563e563e663e163dc63f364013400b3e163df63dd63db63db63da63da63d963d863d763d963dd63e163e763f063f763ff63ee63cc53dd63e763e663e663e563e663e863e863dd63e96400b401b3ff6;
   
   
    fd = $fopen("C:/Users/Asrith S/OneDrive/Desktop/MiniProj/layer1.txt", "r");
    for (i=0; i<6; i=i+1) begin
       code = $fscanf(fd, "%h", memory1[i]);
    end
    for (i = 0; i < 6; i = i + 1) begin
            Conv1F[i*5*5*16+:5*5*16] = memory1[i];
    end

    fd = $fopen("C:/Users/Asrith S/OneDrive/Desktop/MiniProj/layer2.txt", "r");
    for (i=0; i<16; i=i+1) begin
       code = $fscanf(fd, "%h", memory2[i]);
    end
    for (i = 0; i < 16; i = i + 1) begin
            Conv2F[i*5*5*16*6+:5*5*16*6] = memory2[i];
    end

  #(PERIOD/2)
  reset = 1'b0;
  #(PERIOD/2)
  #((7*1457+6*784*6+8+18*22*152 + 6*1600 + 20 + 10000)*PERIOD)
  #(PERIOD*1204) 
  $stop;
  
end

Lenet UUT 
(
	.clk(clk),
	.reset(reset),
	.CNNinput(input_ANN),
	.Conv1F(Conv1F),
	.Conv2F(Conv2F),
	.LeNetoutput(output_ANN)
);

endmodule 